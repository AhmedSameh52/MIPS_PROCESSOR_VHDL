library IEEE;
use IEEE.STD_LOGIC_1164.ALL;


entity Decoder1 is
    Port ( Input : in  STD_LOGIC_VECTOR (4 downto 0);
           E : in  STD_LOGIC;
           O : out  STD_LOGIC_VECTOR (31 downto 0));
end Decoder1;

architecture Behavioral of Decoder1 is

begin

O <= (others=> 'Z') WHEN E = '0'
ELSE
"00000000000000000000000000000001" WHEN Input = "00000" ELSE
"00000000000000000000000000000010" WHEN Input = "00001" ELSE
"00000000000000000000000000000100" WHEN Input = "00010" ELSE
"00000000000000000000000000001000" WHEN Input = "00011" ELSE
"00000000000000000000000000010000" WHEN Input = "00100" ELSE
"00000000000000000000000000100000" WHEN Input = "00101" ELSE
"00000000000000000000000001000000" WHEN Input = "00110" ELSE
"00000000000000000000000010000000" WHEN Input = "00111" ELSE
"00000000000000000000000100000000" WHEN Input = "01000" ELSE
"00000000000000000000001000000000" WHEN Input = "01001" ELSE
"00000000000000000000010000000000" WHEN Input = "01010" ELSE
"00000000000000000000100000000000" WHEN Input = "01011" ELSE
"00000000000000000001000000000000" WHEN Input = "01100" ELSE
"00000000000000000010000000000000" WHEN Input = "01101" ELSE
"00000000000000000100000000000000" WHEN Input = "01110" ELSE
"00000000000000001000000000000000" WHEN Input = "01111" ELSE
"00000000000000010000000000000000" WHEN Input = "10000" ELSE
"00000000000000100000000000000000" WHEN Input = "10001" ELSE
"00000000000001000000000000000000" WHEN Input = "10010" ELSE
"00000000000010000000000000000000" WHEN Input = "10011" ELSE
"00000000000100000000000000000000" WHEN Input = "10100" ELSE
"00000000001000000000000000000000" WHEN Input = "10101" ELSE
"00000000010000000000000000000000" WHEN Input = "10110" ELSE
"00000000100000000000000000000000" WHEN Input = "10111" ELSE
"00000001000000000000000000000000" WHEN Input = "11000" ELSE
"00000010000000000000000000000000" WHEN Input = "11001" ELSE
"00000100000000000000000000000000" WHEN Input = "11010" ELSE
"00001000000000000000000000000000" WHEN Input = "11011" ELSE
"00010000000000000000000000000000" WHEN Input = "11100" ELSE
"00100000000000000000000000000000" WHEN Input = "11101" ELSE
"01000000000000000000000000000000" WHEN Input = "11110" ELSE
"10000000000000000000000000000000" WHEN Input = "11111" ELSE

(others => 'Z');

end Behavioral;